* C:\FOSSEE\eSim\library\SubcircuitLibrary\xor_gate\xor_gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 2/2/2022 10:50:46 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M14-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M14-Pad1_ mosfet_p		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND mosfet_n		
M4  Net-_M14-Pad1_ Net-_M3-Pad2_ Net-_M11-Pad2_ Net-_M14-Pad1_ mosfet_p		
M3  Net-_M11-Pad2_ Net-_M3-Pad2_ GND GND mosfet_n		
M14  Net-_M14-Pad1_ Net-_M10-Pad3_ Net-_M13-Pad1_ Net-_M14-Pad1_ mosfet_p		
M13  Net-_M13-Pad1_ Net-_M10-Pad3_ GND GND mosfet_n		
M7  Net-_M14-Pad1_ Net-_M3-Pad2_ Net-_M10-Pad1_ Net-_M14-Pad1_ mosfet_p		
M8  Net-_M10-Pad1_ Net-_M11-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad1_ mosfet_p		
M9  Net-_M14-Pad1_ Net-_M1-Pad1_ Net-_M10-Pad1_ Net-_M14-Pad1_ mosfet_p		
M10  Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad1_ mosfet_p		
M5  Net-_M10-Pad3_ Net-_M3-Pad2_ Net-_M5-Pad3_ Net-_M5-Pad3_ mosfet_n		
M6  Net-_M5-Pad3_ Net-_M1-Pad1_ GND GND mosfet_n		
M11  Net-_M10-Pad3_ Net-_M11-Pad2_ Net-_M11-Pad3_ Net-_M11-Pad3_ mosfet_n		
M12  Net-_M11-Pad3_ Net-_M1-Pad2_ GND GND mosfet_n		
U1  Net-_M1-Pad2_ Net-_M3-Pad2_ Net-_M13-Pad1_ PORT		
v1  Net-_M14-Pad1_ GND 3.3v		

.end
